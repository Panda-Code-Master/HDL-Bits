module top_module( 
    input wire a,b,c,
    output reg w,x,y,z );
  
    assign w = a ;
    assign x = b ;
    assign y = b ;
    assign z = c ;
           
endmodule
